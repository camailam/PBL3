module seven_segment_decoder (
    input [3:0] input_number,  // 4-bit input representing numbers 0 to 9
    output reg [6:0] seg_display // 7-bit output for controlling seven-segment display
);

always @* begin
    case(input_number)
        4'b0000: seg_display = 7'b1000000; // 0
        4'b0001: seg_display = 7'b1111001; // 1
        4'b0010: seg_display = 7'b0100100; // 2
        4'b0011: seg_display = 7'b0110000; // 3
        4'b0100: seg_display = 7'b0011001; // 4
        4'b0101: seg_display = 7'b0010010; // 5
        4'b0110: seg_display = 7'b0000010; // 6
        4'b0111: seg_display = 7'b1111000; // 7
        4'b1000: seg_display = 7'b0000000; // 8
        4'b1001: seg_display = 7'b0010000; // 9
        default: seg_display = 7'b1111111;  // Invalid input
    endcase
end

endmodule 